* ============================================================================
* RETIFICADORES - Meia Onda, Onda Completa e Ponte Retificadora
* ============================================================================
*
* DESCRICAO:
* ----------
* Este circuito demonstra os três tipos principais de retificadores usados
* em fontes de alimentação para converter AC em DC. Compara desempenho,
* ripple e eficiência de cada topologia.
*
* TOPOLOGIAS:
* -----------
* 1. RETIFICADOR MEIA ONDA (Half-Wave):
*    - 1 diodo
*    - Conduz apenas no semiciclo positivo
*    - Ripple alto (~121% sem filtro)
*    - Frequência de ripple = frede
*    - Eficiência: ~40.6%
*
* 2. RETIFICADOR PONTE (Bridge Rectifier):
*    - 4 diodos em configuração ponte
*    - Usa ambos os semiciclos
*    - Não precisa de center tap
*    - Ripple médio (~48% sem filtro)
*    - Frequência de ripple = 2 × frede
*    - Eficiência: ~81.2%
*    - Queda de tensão: 2 × Vd (dois diodos em série)
*
* NOTA: Retificador onda completa center-tap removido para evitar problemas
*       de convergência (loop de fontes de tensão). O retificador ponte é
*       funcionalmente equivalente e mais comum na prática.
*
* FILTRO CAPACITIVO:
* ------------------
* Adiciona capacitor na saída para suavizar o ripple:
*   - Ripple reduzido para ~1-10% (dependendo de C e Iload)
*   - Ripple voltage: Vr ≈ Iload / (f × C)
*   - Fator de ripple: r = Vr / Vdc
*
* PARAMETROS IMPORTANTES:
* -----------------------
*   - PIV (Peak Inverse Voltage): tensão reversa máxima no diodo
*   - Ripple factor: relação entre AC e DC na saída
*   - Regulation: variação de Vout com a carga
*
* AUTOR: Leonardo Araujo
* DATA: 2025-12-17
* ============================================================================

.title Retificadores - Meia Onda, Onda Completa e Ponte

* ============================================================================
* OPCOES DE SIMULACAO
* ============================================================================
* Opções melhoradas para convergência com retificadores
.options POST RELTOL=1e-3 ABSTOL=1e-9 VNTOL=1e-4
.options TRTOL=7 ITL1=300 ITL2=200 ITL4=100

* ============================================================================
* FONTE AC (Rede Elétrica - 60Hz, 12Vrms ≈ 17Vpk)
* ============================================================================
* Simula secundário de transformador 12V AC
VAC_HW ac_hw 0 SIN(0 17 60 0 0)      ; Para meia onda
VAC_BR ac_br 0 SIN(0 17 60 0 0)      ; Para ponte

* ============================================================================
* RETIFICADOR MEIA ONDA (SEM FILTRO)
* ============================================================================
* Topologia: AC --[D1]--> out --[Rload]--> GND

D_HW ac_hw out_hw DMOD
Rload_HW out_hw 0 1k

* ============================================================================
* RETIFICADOR MEIA ONDA (COM FILTRO CAPACITIVO)
* ============================================================================
* Filtro: capacitor de 470uF + resistência de bleed

D_HWF ac_hw out_hwf DMOD
Cfilt_HWF out_hwf 0 470u
Rbleed_HWF out_hwf 0 100k    ; Resistência de bleed para convergência
Rload_HWF out_hwf 0 1k

* ============================================================================
* RETIFICADOR PONTE (SEM FILTRO)
* ============================================================================
* Topologia correta de ponte retificadora:
*   D1: AC → top_node
*   D2: GND → top_node
*   D3: bot_node → AC
*   D4: bot_node → GND
*   Carga: entre top_node e bot_node

D_BR1 ac_br n_br_top DMOD     ; AC → nó superior
D_BR2 0 n_br_top DMOD         ; GND → nó superior
D_BR3 n_br_bot ac_br DMOD     ; nó inferior → AC
D_BR4 n_br_bot 0 DMOD         ; nó inferior → GND
Rload_BR n_br_top n_br_bot 1k ; Carga entre top e bottom
Rgnd_BR n_br_bot 0 1Meg       ; Referência ao GND (alta impedância)

* ============================================================================
* RETIFICADOR PONTE (COM FILTRO)
* ============================================================================

D_BRF1 ac_br n_brf_top DMOD
D_BRF2 0 n_brf_top DMOD
D_BRF3 n_brf_bot ac_br DMOD
D_BRF4 n_brf_bot 0 DMOD
Cfilt_BRF n_brf_top n_brf_bot 470u  ; Filtro entre top e bottom
Rload_BRF n_brf_top n_brf_bot 1k
Rgnd_BRF n_brf_bot 0 1Meg             ; Referência ao GND

* ============================================================================
* MODELO DO DIODO
* ============================================================================
* Diodo de silício genérico (1N4007-like)
.model DMOD D(
+ IS=1e-14      ; Corrente de saturação
+ RS=0.05       ; Resistência série (Ohms)
+ N=1.7         ; Coeficiente de emissão
+ BV=1000       ; Tensão de breakdown (V)
+ IBV=1e-3      ; Corrente de breakdown (A)
+ VJ=0.7        ; Tensão de junção (V)
+ CJO=15p       ; Capacitância de junção (F)
+ TT=5n         ; Tempo de trânsito (s)
+ )

* ============================================================================
* ANALISE TRANSIENTE
* ============================================================================
* Simular 5 ciclos (5/60Hz = 83.3ms)
* Timestep inicial: 10us, tempo total: 83.3ms, timestep máximo: 100us
.tran 10u 83.3m 0 100u

* ============================================================================
* MEDICOES
* ============================================================================
* Valores médios (DC) e ripple

.measure tran Vdc_hw AVG v(out_hw) FROM=33.3m TO=83.3m
.measure tran Vdc_hwf AVG v(out_hwf) FROM=33.3m TO=83.3m
.measure tran Vdc_br AVG v(n_br_top) FROM=33.3m TO=83.3m
.measure tran Vdc_brf AVG v(n_brf_top) FROM=33.3m TO=83.3m

* Ripple (pico a pico)
.measure tran Vripple_hw PP v(out_hw) FROM=33.3m TO=83.3m
.measure tran Vripple_hwf PP v(out_hwf) FROM=33.3m TO=83.3m
.measure tran Vripple_br PP v(n_br_top) FROM=33.3m TO=83.3m
.measure tran Vripple_brf PP v(n_brf_top) FROM=33.3m TO=83.3m

* ============================================================================
* PLOTS E ANALISE
* ============================================================================
.control
run

* Plot 1: Entrada AC
plot v(ac_hw)
+ title "Entrada AC - 12Vrms (17Vpk) @ 60Hz" xlabel "Tempo (ms)" ylabel "Tensao (V)"

* Plot 2: Comparação Meia Onda (sem e com filtro)
plot v(out_hw) v(out_hwf)
+ title "Retificador Meia Onda - Sem Filtro vs Com Filtro 470uF" xlabel "Tempo (ms)" ylabel "Tensao (V)"

* Plot 3: Comparação Ponte (sem e com filtro)
plot v(n_br_top,n_br_bot) v(n_brf_top,n_brf_bot)
+ title "Retificador Ponte - Sem Filtro vs Com Filtro 470uF" xlabel "Tempo (ms)" ylabel "Tensao (V)"

* Plot 4: Comparação de todas as topologias COM filtro
plot v(out_hwf) v(n_brf_top,n_brf_bot)
+ title "Comparacao: Meia Onda vs Ponte (com filtro)" xlabel "Tempo (ms)" ylabel "Tensao (V)"

* Plot 5: Zoom no ripple (últimos 2 ciclos)
plot v(out_hwf) v(n_brf_top,n_brf_bot) xlimit 50m 83.3m
+ title "Ripple - Zoom nos ultimos 2 ciclos" xlabel "Tempo (ms)" ylabel "Tensao (V)"

* Exportar dados para CSV
set wr_singlescale
set wr_vecnames
option numdgt=7
wrdata circuits/09_fontes_alimentacao/retificadores_saidas.csv v(out_hw) v(out_hwf) v(n_br_top,n_br_bot) v(n_brf_top,n_brf_bot)
wrdata circuits/09_fontes_alimentacao/retificadores_entrada.csv v(ac_hw)

echo ""
echo "============================================================================"
echo "RESULTADOS DOS RETIFICADORES"
echo "============================================================================"
echo ""
echo "RETIFICADOR MEIA ONDA:"
echo "  Sem filtro - Vdc:" Vdc_hw "V, Ripple:" Vripple_hw "V"
echo "  Com filtro - Vdc:" Vdc_hwf "V, Ripple:" Vripple_hwf "V"
echo ""
echo "RETIFICADOR PONTE:"
echo "  Sem filtro - Vdc:" Vdc_br "V, Ripple:" Vripple_br "V"
echo "  Com filtro - Vdc:" Vdc_brf "V, Ripple:" Vripple_brf "V"
echo ""
echo "OBSERVACOES:"
echo "  - Meia onda: ripple @ 60Hz (frede)"
echo "  - Ponte: ripple @ 120Hz (2×frede)"
echo "  - Filtro capacitivo reduz ripple significativamente"
echo "  - Ponte: 2 diodos em serie = maior queda de tensao (~1.4V)"
echo "============================================================================"
echo ""

print Vdc_hw Vdc_hwf Vdc_br Vdc_brf

quit
.endc

.end
