"RC Low-Pass Filter"
* Simple RC network

V1 in 0 1
R1 in out 1k
C1 out 0 1u

.end
