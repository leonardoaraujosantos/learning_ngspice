* ==============================================================
* RLC TRANSIENTE (RINGING) — “não é oscilador”, é oscilação amortecida
* Objetivo:
*   1) Aplicar um degrau de 0V -> 10V (simula “ligar” a fonte DC)
*   2) Observar a oscilação natural do circuito RLC e seu decaimento
*   3) Rodar por ~10 ciclos (≈ 31.4 s) e medir tensão em 2 instantes:
*        - depois de ~10 ciclos (31.4 s)
*        - no final da simulação (35 s)
*
* Circuito:
*   V1 (degrau) -> L1 (série) -> nó OUT
*   nó OUT ligado a R1 || C1 para o GND
* ==============================================================

* ---------- Fonte ----------
* PWL cria um degrau: em t=0 está 0V e em t=1us sobe para 10V.
* Isso evita o SPICE iniciar direto em regime estacionário.
V1 in 0 PWL(0 0 1u 10)

* ---------- Indutor em série ----------
* 500 mH = 0.5 H
L1 in out 500m

* ---------- Carga no nó OUT ----------
* Capacitor para o terra (500 mF = 0.5 F)
C1 out 0 500m

* Resistor para o terra (10 Ω) — fornece amortecimento (dissipa energia)
* Valor reduzido de 10k para 10 para aumentar amortecimento (zeta ≈ 0.1)
R1 out 0 10

* ---------- Análise Transiente ----------
* Passo de amostragem (TSTEP) = 1 ms (obrigatoriamente > 0 no NGspice)
* Tempo final = 15 s (≈ 5 ciclos completos, porque T ≈ 3.14 s)
.tran 1m 15

* ---------- Cálculo de referência ----------
* Frequência natural aproximada:
*   f0 = 1 / (2*pi*sqrt(L*C))
*   L=0.5 H, C=0.5 F  => f0 ≈ 0.318 Hz
* Período aproximado:
*   T ≈ 1/f0 ≈ 3.14 s
* 10 ciclos => ~31.4 s
*
* (A presença de R muda um pouco a frequência amortecida, mas é próximo.)

* ---------- Medições (.measure) ----------
* Mede picos para visualizar o decaimento do envelope:

* Primeiro pico (1º ciclo):
.measure tran Vout_peak_1st MAX v(out) FROM=0 TO=3.14

* Tensão RMS no 1º ciclo:
.measure tran Vout_RMS_1st RMS v(out) FROM=0 TO=3.14

* Depois de 2 ciclos (~6.28s):
.measure tran Vout_after_2cycles FIND v(out) AT=6.28

* Pico após 2 ciclos (3º ciclo):
.measure tran Vout_peak_3rd MAX v(out) FROM=6.28 TO=9.42

* Tensão RMS no 3º ciclo:
.measure tran Vout_RMS_3rd RMS v(out) FROM=6.28 TO=9.42

* Depois de 4 ciclos (~12.56s):
.measure tran Vout_after_4cycles FIND v(out) AT=12.56

* Tensão RMS no período final (últimos 3s):
.measure tran Vout_RMS_final RMS v(out) FROM=12 TO=15

* Tensão no final da simulação:
.measure tran Vout_end FIND v(out) AT=15

* ---------- Bloco de controle (para rodar, plotar e salvar) ----------
.control
  run

  * Se você rodar em modo interativo (ngspice arquivo.cir),
  * este comando abre/mostra o gráfico:
  plot v(out)

  * Salva dados em arquivo para plotar fora (gnuplot/python):
  wrdata vout.dat time v(out)

  * Mostra na tela (útil no modo interativo; no batch as .measure já aparecem):
  echo "==== DECAIMENTO DA OSCILAÇÃO ===="
  echo ""
  echo "1º CICLO:"
  echo "  Pico              = " Vout_peak_1st
  echo "  RMS               = " Vout_RMS_1st
  echo ""
  echo "APÓS 2 CICLOS (6.28s):"
  echo "  V(out)            = " Vout_after_2cycles
  echo ""
  echo "3º CICLO:"
  echo "  Pico              = " Vout_peak_3rd
  echo "  RMS               = " Vout_RMS_3rd
  echo ""
  echo "APÓS 4 CICLOS (12.56s):"
  echo "  V(out)            = " Vout_after_4cycles
  echo ""
  echo "PERÍODO FINAL (12-15s):"
  echo "  RMS               = " Vout_RMS_final
  echo "  V(out) em t=15s   = " Vout_end
.endc

.end
