* ============================================================================
* Teste de Diodo Simples usando Verilog-A
* ============================================================================
*
* COMPILAR:
*   openvaf diodo_simples.va
*
* EXECUTAR:
*   ngspice teste_diodo.cir
*
* ============================================================================

.title Teste de Diodo Verilog-A

* Carregar modelo compilado
.pre_osdi diodo_simples.osdi

* Retificador de meia onda
Vin in 0 SIN(0 5 60)
D1 in out diodo_simples Is=1e-14 n=1.0 Rs=10 Cj0=10p
Rload out 0 1k
Cfilt out 0 100u

* Analises
.tran 1m 50m
.dc Vin -1 1 0.01

.control
  * Analise transiente
  tran 1m 50m
  set curplot = tran1

  plot v(in) v(out) title 'Retificador de Meia Onda'
  plot i(Vin) title 'Corrente no Diodo'

  * Medicoes transiente
  meas tran Vpico_in MAX v(in)
  meas tran Vpico_out MAX v(out)
  meas tran Vripple PP v(out) FROM=33.3m TO=50m

  echo "======================================"
  echo "Analise Transiente - Retificador"
  echo "======================================"
  echo "Tensao de pico entrada: " $&Vpico_in " V"
  echo "Tensao de pico saida:   " $&Vpico_out " V"
  echo "Ripple:                 " $&Vripple " V"

  * Analise DC - Curva I-V
  dc Vin -1 1 0.01
  set curplot = dc1

  plot i(Vin) vs v(in) title 'Curva I-V do Diodo' xlabel 'Tensao (V)' ylabel 'Corrente (A)'

  * Escala logaritmica para ver corrente reversa
  let I_abs = abs(i(Vin))
  plot I_abs vs v(in) ylog title 'Curva I-V (log)' xlabel 'Tensao (V)' ylabel 'Corrente (A)'

  * Exportar dados
  wrdata diodo_iv.csv v(in) i(Vin)

  * Medicoes DC
  meas dc I_forward find i(Vin) at=0.7
  meas dc I_reverse find i(Vin) at=-1

  echo "======================================"
  echo "Analise DC - Curva I-V"
  echo "======================================"
  echo "Corrente em +0.7V: " $&I_forward " A"
  echo "Corrente em -1.0V: " $&I_reverse " A"
.endc

.end
