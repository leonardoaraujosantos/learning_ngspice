* Filtro RC Passa-Baixa - Esquematico Simples
* Vin -> R -> Vout -> C -> GND

V1 in 0 DC 1 AC 1
R1 in out 1k
C1 out 0 100n

.end
