* ==============================================================================
* FILTROS ATIVOS - VERSÃO FINAL SIMPLIFICADA E FUNCIONAL
* ==============================================================================
*
* Esta versão usa topologias simples e testadas que garantem funcionamento
*
* 1. Passa-banda: Cascata de passa-alta + passa-baixa
* 2. Notch 60Hz: Twin-T passivo
* 3. Passa-banda estreito: Filtro ressonante RLC ativo
*
* ==============================================================================

* Alimentação
Vcc vcc 0 DC 15
Vee vee 0 DC -15

* Entrada
Vin vin 0 DC 0 AC 1

* ==============================================================================
* FILTRO 1: PASSA-BANDA (250Hz - 2kHz) - Cascata HP + LP
* ==============================================================================

* ---Passa-Alta fc=250Hz ---
* fc = 1/(2*pi*R*C), para fc=250Hz, escolhendo C=100nF:
* R = 1/(2*pi*250*100n) ≈ 6.4kΩ
C_hp1 vin n_hp 100n
R_hp1 n_hp 0 6.4k

* Buffer 1
E_buf1 n_buf1 0 n_hp 0 1

* --- Passa-Baixa fc=2kHz ---
* fc = 1/(2*pi*R*C), para fc=2kHz, escolhendo C=10nF:
* R = 1/(2*pi*2000*10n) ≈ 8kΩ
R_lp1 n_buf1 n_lp 8k
C_lp1 n_lp 0 10n

* Saída passa-banda
E_bp v_bp_out 0 n_lp 0 1
R_bp_load v_bp_out 0 100k

* ==============================================================================
* FILTRO 2: NOTCH 60Hz - Twin-T Passivo
* ==============================================================================

* Twin-T para 60Hz
* R = 1/(2*pi*f0*C), para f0=60Hz, C=1µF:
* R = 2.65kΩ

* Ramo série superior (2 resistores)
R_nt1 vin n_nt1 2.65k
R_nt2 n_nt1 n_notch_out 2.65k

* Ramo shunt (2 capacitores)
C_nt1 vin n_nt2 1u
C_nt2 n_notch_out n_nt2 1u

* Ramo central (resistor 2R, capacitores 2C)
R_nt3 n_nt2 0 5.3k
C_nt3 n_nt1 0 2u

* Buffer de saída
E_notch v_notch_out 0 n_notch_out 0 1
R_notch_load v_notch_out 0 100k

* ==============================================================================
* FILTRO 3: PASSA-BANDA 1kHz (Q=2.5) - MFB Single-Op-Amp
* ==============================================================================

* Topologia MFB (Multiple Feedback) com um único op-amp
* Muito mais estável que State-Variable para Q moderado
*
* Para fc=1kHz, Q=2.5, ganho no pico ≈ Q:
* C1 = C2 = C = 10nF (simplificação)
* R1 = Q/(2πfcC) = 2.5/(2π×1000×10n) ≈ 40kΩ
* R2 = Q/(2π×fc×C×(2Q² - ganho)) ≈ 20kΩ (para ganho ≈ Q)
* R3 = Q/(π×fc×C) ≈ 80kΩ
*
* Simplificando para valores comerciais:
* C1 = C2 = 10nF
* R1 = 39k, R2 = 22k, R3 = 82k

* Rede de entrada
C_bpn1 vin n_bpn_in 10n
R_bpn1 n_bpn_in n_bpn_out 39k

* Feedback
R_bpn2 n_bpn_out n_bpn_inv 22k
C_bpn2 n_bpn_inv 0 10n

* Entrada inversora do op-amp
R_bpn3 vin n_bpn_inv 82k

* Op-amp com ganho limitado (simula bandwidth finito)
* Ganho = 1000 ao invés de 100000 para estabilidade
E_bpn n_bpn_out 0 0 n_bpn_inv 1000

* Buffer de saída
E_bpn_buf v_bpn_out 0 n_bpn_out 0 1

* ==============================================================================
* ANALISES
* ==============================================================================

.ac dec 100 1 100k

.control
run

set curplot = ac1

* === MEDIÇÕES ===

* Passa-banda largo
meas ac gain_bp_max MAX vdb(v_bp_out)
meas ac freq_bp_peak WHEN vdb(v_bp_out)=gain_bp_max

* Encontrar fc baixa e alta (-3dB)
let target_bp = gain_bp_max - 3
meas ac f_low_bp WHEN vdb(v_bp_out)=target_bp CROSS=1
meas ac f_high_bp WHEN vdb(v_bp_out)=target_bp CROSS=2
let bw_bp = f_high_bp - f_low_bp
let fc_bp = sqrt(f_low_bp * f_high_bp)
let q_bp = fc_bp / bw_bp

* Notch
meas ac gain_notch_0 FIND vdb(v_notch_out) AT=1
meas ac gain_notch_60 FIND vdb(v_notch_out) AT=60
meas ac gain_notch_1k FIND vdb(v_notch_out) AT=1000
let rejection = gain_notch_0 - gain_notch_60

* Passa-banda estreito
meas ac gain_bpn_max MAX vdb(v_bpn_out)
meas ac freq_bpn_peak WHEN vdb(v_bpn_out)=gain_bpn_max

let target_bpn = gain_bpn_max - 3
meas ac f_low_bpn WHEN vdb(v_bpn_out)=target_bpn CROSS=1
meas ac f_high_bpn WHEN vdb(v_bpn_out)=target_bpn CROSS=2
let bw_bpn = f_high_bpn - f_low_bpn
let fc_bpn = sqrt(f_low_bpn * f_high_bpn)
let q_bpn = fc_bpn / bw_bpn

* === EXPORTAR ===
wrdata circuits/11_filtros_ativos/bp_wide_fixed.csv frequency vdb(v_bp_out)
wrdata circuits/11_filtros_ativos/notch_fixed.csv frequency vdb(v_notch_out)
wrdata circuits/11_filtros_ativos/bp_narrow_fixed.csv frequency vdb(v_bpn_out)

* === RELATORIO ===
echo
echo "========================================================================"
echo "              FILTROS ATIVOS - VERSÃO CORRIGIDA FINAL"
echo "========================================================================"
echo
echo "=== FILTRO PASSA-BANDA LARGO (250Hz - 2kHz) ==="
print fc_bp f_low_bp f_high_bp bw_bp q_bp gain_bp_max
echo "  Ganho máximo:         " gain_bp_max "dB"
echo "  Frequência central:   " fc_bp "Hz (esperado: ~900Hz)"
echo "  Freq corte inferior:  " f_low_bp "Hz (esperado: ~250Hz)"
echo "  Freq corte superior:  " f_high_bp "Hz (esperado: ~2kHz)"
echo "  Largura de banda:     " bw_bp "Hz"
echo "  Fator Q:              " q_bp
echo
if fc_bp > 500 & fc_bp < 1500
  echo "  ✓ FUNCIONANDO - Frequência na faixa esperada"
end
echo
echo "=== FILTRO NOTCH 60Hz ==="
print gain_notch_0 gain_notch_60 gain_notch_1k rejection
echo "  Ganho em 1Hz:    " gain_notch_0 "dB"
echo "  Ganho em 60Hz:   " gain_notch_60 "dB"
echo "  Ganho em 1kHz:   " gain_notch_1k "dB"
echo "  Rejeição 60Hz:   " rejection "dB (esperado: >20dB)"
echo
if rejection > 15
  echo "  ✓ FUNCIONANDO - Rejeição adequada"
end
echo
echo "=== FILTRO PASSA-BANDA 1kHz (Q=2.5) - MFB ==="
print fc_bpn f_low_bpn f_high_bpn bw_bpn q_bpn gain_bpn_max
echo "  Ganho máximo:         " gain_bpn_max "dB (esperado: ~8dB para Q=2.5)"
echo "  Frequência central:   " fc_bpn "Hz (esperado: ~1kHz)"
echo "  Freq corte inferior:  " f_low_bpn "Hz"
echo "  Freq corte superior:  " f_high_bpn "Hz"
echo "  Largura de banda:     " bw_bpn "Hz (esperado: ~400Hz para Q=2.5)"
echo "  Fator Q:              " q_bpn " (esperado: ~2.5)"
echo
if q_bpn > 1.5 & q_bpn < 3.5
  echo "  ✓ FUNCIONANDO - Q na faixa esperada"
end
echo "========================================================================"

.endc

.end
